//modulo de saida do processador
module saida (clk,dado,controle,d0,d1,d2,d3,d4,d5,d6,d7,neg);

input clk; //clock do processador
input [31:0]dado; //dado para impressao
input controle; //sinal de controle do modulo de saida
output reg [6:0] d0,d1,d2,d3,d4,d5,d6,d7; //vetores correspondentes aos displays de 7 segmentos
output reg neg; //sinal de valor negativo
reg [31:0] entrada; //dado final para a impressao

initial
begin
	entrada = 32'd0; //inicia imprimindo 0
	neg = 1'd0; //sinal de valor negativ apagado
end

always @(posedge clk) //na borda de subida do clock
begin
	if(controle==1) //eh para imprimir?
	begin
		if(dado[31]==1) //o bit mais significado eh 1? valor negativo
			begin
				entrada = ~(dado-32'd1);
				neg = 1;
			end
		else
			begin //valor positivo
				entrada = dado;
				neg = 0;
			end
	end
end

always@(entrada) // se entrada mudar os displays mudam
	begin
		case (entrada[3:0])
			4'b0000: d0=7'b1000000;
			4'b0001: d0=7'b1111001;
			4'b0010: d0=7'b0100100;
			4'b0011: d0=7'b0110000;
			4'b0100: d0=7'b0011001;
			4'b0101: d0=7'b0010010;
			4'b0110: d0=7'b0000010;
			4'b0111: d0=7'b1111000;
			4'b1000: d0=7'b0000000;
			4'b1001: d0=7'b0010000;
			4'b1010: d0=7'b0001000;
			4'b1011: d0=7'b0000011;
			4'b1100: d0=7'b1000110;
			4'b1101: d0=7'b0100001;
			4'b1110: d0=7'b0000110;
			4'b1111: d0=7'b0001110;
		endcase
		case (entrada[7:4])
			4'b0000: d1=7'b1000000;
			4'b0001: d1=7'b1111001;
			4'b0010: d1=7'b0100100;
			4'b0011: d1=7'b0110000;
			4'b0100: d1=7'b0011001;
			4'b0101: d1=7'b0010010;
			4'b0110: d1=7'b0000010;
			4'b0111: d1=7'b1111000;
			4'b1000: d1=7'b0000000;
			4'b1001: d1=7'b0010000;
			4'b1010: d1=7'b0001000;
			4'b1011: d1=7'b0000011;
			4'b1100: d1=7'b1000110;
			4'b1101: d1=7'b0100001;
			4'b1110: d1=7'b0000110;
			4'b1111: d1=7'b0001110;
		endcase
		case (entrada[11:8])
			4'b0000: d2=7'b1000000;
			4'b0001: d2=7'b1111001;
			4'b0010: d2=7'b0100100;
			4'b0011: d2=7'b0110000;
			4'b0100: d2=7'b0011001;
			4'b0101: d2=7'b0010010;
			4'b0110: d2=7'b0000010;
			4'b0111: d2=7'b1111000;
			4'b1000: d2=7'b0000000;
			4'b1001: d2=7'b0010000;
			4'b1010: d2=7'b0001000;
			4'b1011: d2=7'b0000011;
			4'b1100: d2=7'b1000110;
			4'b1101: d2=7'b0100001;
			4'b1110: d2=7'b0000110;
			4'b1111: d2=7'b0001110;
		endcase
		case (entrada[15:12])
			4'b0000: d3=7'b1000000;
			4'b0001: d3=7'b1111001;
			4'b0010: d3=7'b0100100;
			4'b0011: d3=7'b0110000;
			4'b0100: d3=7'b0011001;
			4'b0101: d3=7'b0010010;
			4'b0110: d3=7'b0000010;
			4'b0111: d3=7'b1111000;
			4'b1000: d3=7'b0000000;
			4'b1001: d3=7'b0010000;
			4'b1010: d3=7'b0001000;
			4'b1011: d3=7'b0000011;
			4'b1100: d3=7'b1000110;
			4'b1101: d3=7'b0100001;
			4'b1110: d3=7'b0000110;
			4'b1111: d3=7'b0001110;
		endcase
		case (entrada[19:16])
			4'b0000: d4=7'b1000000;
			4'b0001: d4=7'b1111001;
			4'b0010: d4=7'b0100100;
			4'b0011: d4=7'b0110000;
			4'b0100: d4=7'b0011001;
			4'b0101: d4=7'b0010010;
			4'b0110: d4=7'b0000010;
			4'b0111: d4=7'b1111000;
			4'b1000: d4=7'b0000000;
			4'b1001: d4=7'b0010000;
			4'b1010: d4=7'b0001000;
			4'b1011: d4=7'b0000011;
			4'b1100: d4=7'b1000110;
			4'b1101: d4=7'b0100001;
			4'b1110: d4=7'b0000110;
			4'b1111: d4=7'b0001110;
		endcase
		case (entrada[23:20])
			4'b0000: d5=7'b1000000;
			4'b0001: d5=7'b1111001;
			4'b0010: d5=7'b0100100;
			4'b0011: d5=7'b0110000;
			4'b0100: d5=7'b0011001;
			4'b0101: d5=7'b0010010;
			4'b0110: d5=7'b0000010;
			4'b0111: d5=7'b1111000;
			4'b1000: d5=7'b0000000;
			4'b1001: d5=7'b0010000;
			4'b1010: d5=7'b0001000;
			4'b1011: d5=7'b0000011;
			4'b1100: d5=7'b1000110;
			4'b1101: d5=7'b0100001;
			4'b1110: d5=7'b0000110;
			4'b1111: d5=7'b0001110;
		endcase
		case (entrada[27:24])
			4'b0000: d6=7'b1000000;
			4'b0001: d6=7'b1111001;
			4'b0010: d6=7'b0100100;
			4'b0011: d6=7'b0110000;
			4'b0100: d6=7'b0011001;
			4'b0101: d6=7'b0010010;
			4'b0110: d6=7'b0000010;
			4'b0111: d6=7'b1111000;
			4'b1000: d6=7'b0000000;
			4'b1001: d6=7'b0010000;
			4'b1010: d6=7'b0001000;
			4'b1011: d6=7'b0000011;
			4'b1100: d6=7'b1000110;
			4'b1101: d6=7'b0100001;
			4'b1110: d6=7'b0000110;
			4'b1111: d6=7'b0001110;
		endcase
		case (entrada[31:28])
			4'b0000: d7=7'b1000000;
			4'b0001: d7=7'b1111001;
			4'b0010: d7=7'b0100100;
			4'b0011: d7=7'b0110000;
			4'b0100: d7=7'b0011001;
			4'b0101: d7=7'b0010010;
			4'b0110: d7=7'b0000010;
			4'b0111: d7=7'b1111000;
			4'b1000: d7=7'b0000000;
			4'b1001: d7=7'b0010000;
			4'b1010: d7=7'b0001000;
			4'b1011: d7=7'b0000011;
			4'b1100: d7=7'b1000110;
			4'b1101: d7=7'b0100001;
			4'b1110: d7=7'b0000110;
			4'b1111: d7=7'b0001110;
		endcase
	end
endmodule